

module IEEE_adder_tb;

    timeunit 1ns/1ps;
    localparam CLK_PERIOD = 10;
    logic command;
    logic clk=0;
    logic [31:0] number1;
    logic [31:0] number2;
    logic [31:0] sum;
    
    IEEE_adder dut(.*);

    initial forever #(CLK_PERIOD/2) clk <= !clk;

    initial begin
        @(posedge clk);
        number1 <= 32'b01000000111100000000000000000000; //1 10000001 11100000000000000000000
        number2 <= 32'b11000000001000000000000000000000; //1 10000000 01000000000000000000000
        command <= 1;
                
        #200;
        
        @(posedge clk);
        number1 <= 32'b01000000111100000000000000000000; //0 10000001 11010000000000000000000
        number2 <= 32'b01000000001000000000000000000000; //1 01111110 01000000000000000000000
        command <= 1;
        
        #100;
        @(posedge clk);
        number1 <= 32'b01000000001000000000000000000000; //0 10000001 11010000000000000000000         01000000111100000000000000000000
        number2 <= 32'b01000000111100000000000000000000; //1 01111110 01000000000000000000000
        command <= 1;
        
//        #100;
//        @(posedge clk);
//        number1 <= 32'b00111111100011001110110110010001; //0 10000001 11010000000000000000000         01000000111100000000000000000000
//        number2 <= 32'b00111111100011001100110011001101; //1 01111110 01000000000000000000000
//        command <= 1;

        #100;
        @(posedge clk);
        number1 <= 32'b00111111100011001100110011001101; //0 10000001 11010000000000000000000         01000000111100000000000000000000
        number2 <= 32'b00111111100011001110110110010001; //1 01111110 01000000000000000000000
        command <= 0;       
        
//        @(posedge clk);
//        number1 <= 32'b00111111100011001110110110010001; //0 10000001 11010000000000000000000
//        number2 <= 32'b00111111100011001100110011001101; //1 01111110 01000000000000000000000
//        command <= 0;



        
    end


    
endmodule