module uart_with_rx_parity #(
  parameter CLOCKS_PER_PULSE = 4, //200_000_000/9600
            BITS_PER_WORD    = 8,
            W_OUT //R*C*W_K + C*W_X,
)(
    input  logic clk, rstn, rx,
    output logic m_valid, parity_bit,
    output logic [W_OUT-1:0] m_data
);
    localparam  NUM_WORDS = W_OUT/BITS_PER_WORD;

  // Counters



  // State Machine

    enum {IDLE, START, DATA, PARITY, END} state;

    logic [$clog2(CLOCKS_PER_PULSE) -1:0] c_clocks;
    logic [$clog2(BITS_PER_WORD)    -1:0] c_bits  ;
    logic [$clog2(NUM_WORDS)        -1:0] c_words ;


    always_ff @(posedge clk or negedge rstn) begin
    
    if (!rstn) begin
        {c_words, c_bits, c_clocks, m_valid, m_data} <= '0;
        state <= IDLE;
    end else begin
        m_valid <= 0;
      
            case (state)

            IDLE :  if (rx == 0)                      
                    state <= START;

            START:  if (c_clocks == CLOCKS_PER_PULSE/2-1) begin
                    state <= DATA;
                    c_clocks <= 0;
                end else
                    c_clocks <= c_clocks + 1;

            DATA :  if (c_clocks == CLOCKS_PER_PULSE-1) begin
                    c_clocks <= 0;
                    m_data   <= {rx, m_data[W_OUT-1:1]};   //shift register to add rx after clock cycles of pulse passes

                    if (c_bits == BITS_PER_WORD-1) begin
                        state  <= PARITY;
                        c_bits <= 0;

                        if (c_words == NUM_WORDS-1) begin
                            m_valid <= 1;
                            c_words <= 0;

                        end else 
                            c_words <= c_words + 1;
                    end else 
                        c_bits <= c_bits + 1;
                end else 
                    c_clocks <= c_clocks + 1;
            
//            PARITY : if (rx == ^m_data[BITS_PER_WORD +: BITS_PER_WORD] & c_clocks == CLOCKS_PER_PULSE - 1) begin   //st this state rx is the parity bit
//                        state <= END;
//                        c_clocks <= 0;
//                    end
//                    else if (^m_data[BITS_PER_WORD +: BITS_PER_WORD] != rx & c_clocks == CLOCKS_PER_PULSE - 1) begin
//                        state <= IDLE;
//                        c_clocks <= 0;
                    
//                    end else
//                        c_clocks <= c_clocks + 1;

             PARITY:
                     if (c_clocks == CLOCKS_PER_PULSE-1) begin
                         c_clocks <= 0;
                         parity_bit = ^m_data[BITS_PER_WORD +: BITS_PER_WORD];
                         if (rx == parity_bit) begin
                             state <= END;
                         end else 
                             state <= IDLE; 
                     end else 
                         c_clocks <= c_clocks + 1;    

                    
            END  :  if (c_clocks == CLOCKS_PER_PULSE-1) begin
                        state <= IDLE;
                        c_clocks <= 0;
                    end else
                        c_clocks <= c_clocks + 1;
            endcase
        end
    end
endmodule