module Adder_8bit (
    input logic
);
    
endmodule